`ifndef __FETCH_DECODE_SV
`define __FETCH_DECODE_SV

`ifdef VERILATOR
`include "include/common.sv"
`include "include/pipes.sv"
`else

`endif

module fetch_decode 
    import common::*;
    import pipes::*;(

    
);
    
endmodule

`endif