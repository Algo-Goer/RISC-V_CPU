`ifndef __PIPES_SV
`define __PIPES_SV

`ifdef VERILATOR
`include "include/common.sv"
`endif
package pipes;
	import common::*;
/* Define instrucion decoding rules here */

// parameter F7_RI = 7'bxxxxxxx;
parameter F7_I_TYPE = 7'b0010011;
parameter F7_R_TYPE = 7'b0110011;
parameter F7_LUI = 7'b0110111;
parameter F7_AUIPC = 7'b0010111;
parameter F7_LD = 7'b0000011;
parameter F7_SD = 7'b0100011;
parameter F7_JAL = 7'b1101111;
parameter F7_JALR = 7'b1100111;
parameter F7_BEQ = 7'b1100011;

parameter F7_ADD = 7'b0000000;
parameter F7_SUB = 7'b0100000;
parameter F3_ADD = 3'b000;
parameter F3_AND = 3'b111;
parameter F3_OR = 3'b110;
parameter F3_XOR = 3'b100;


/* Define pipeline structures here */
// alu进行的操作类型
typedef enum logic [4:0] {
	ALU_ADD, ALU_SUB, 
	ALU_OR, ALU_AND, ALU_XOR,
	ALU_EQUAL
} alufunc_t;

// decode判断出的指令类型
typedef enum logic [5 : 0] { 
	UNKNOWN, 
	ADDI, ORI, ANDI, XORI, 
	LUI, AUIPC,
	ADD, SUB, OR, AND, XOR,
	LD, SD,
	JAL, JALR, 
	BEQ
} decode_op_t;

// decode流水段产生的控制信号
typedef struct packed {
    // 指令信息
    decode_op_t op;
    // fetch控制信号
    u1 jump;					//无条件跳转
    // execute控制信号
    alufunc_t func;				// alu操作
    u1 srca_r; 
    u1 srcb_r;                  //两个操作数是否可能需要更新
    // memory控制信号
    u1 memread;					// 内存读使能
    u1 memwrite;				// 内存写使能
    // writeback控制信号
    u1 regwrite;				// regfile写使能
    creg_addr_t dst;			// 写回regfile编号
} decode_control_t;

// execute阶段传递的控制信号
typedef struct packed {
    // fetch控制信号
    u1 jump;					// 条件跳转
    // memory控制信号
    u1 memread;					// 内存读使能
    u1 memwrite;				// 内存写使能
    // writeback控制信号
    u1 regwrite;				// regfile写使能
    creg_addr_t dst;			// 写回regfile编号
} execute_control_t;

// fetch阶段产生的信号
typedef struct packed {
	u32 instruction;			//指令
	u64 pc;						//pc
} fetch_data_t;

// decode阶段产生的信号
typedef struct packed {
    u32 pc;
	creg_addr_t ra1;
    creg_addr_t ra2;
    word_t srca, srcb;			// 操作数
    word_t imm;                 //立即数扩展结果
    word_t pcdata;              // 待计算pc的数据，x[instruction[19 : 15]]
    word_t memdata;				// 待写入内存的数据，x[instruction[24 : 20]]
    decode_control_t ctl;		// 控制信号
} decode_data_t;

// execute阶段产生的信号
typedef struct packed {
    u64 j_addr;                 //跳转地址
    word_t memdata;				// 待写入内存的数据
    word_t result;				// 计算结果，可能作为访存地址，也可能作为regfile写回数据
    execute_control_t ctl;		// 控制信号
} execute_data_t;

// memory阶段产生的信号
typedef struct packed {
	u1 regwrite;				// regfile写使能
	creg_addr_t dst;			// 写回regfile编号
	word_t regdata;				// 写回的数据
	// word_t memdata;				// 待写入内存的数据
} memory_data_t;

// writeback阶段产生的信号
typedef struct packed {
	u1 regwrite;				// regfile写使能
	creg_addr_t dst;			// 写回regfile编号
	word_t regdata;				// 写回的数据
	// word_t memdata;				// 待写入内存的数据
} writeback_data_t;

// forward寄存器模块输入
typedef struct packed {
    u1 valid;
    creg_addr_t dst;
    word_t data;
} forward_data_out;

// hazard寄存器模块输入输出
typedef struct packed {
    creg_addr_t rs, rt;
    creg_addr_t dst;
    u1 regwrite;
    u1 memread;
    u1 jump;
} hazard_data_in;

typedef struct packed {
    u1 stall;
    u1 clear1;
    u1 clear2;
    u1 srca_mux;
    word_t srca_forward;
    u1 srcb_mux;
    word_t srcb_forward;
} hazard_data_out;

endpackage

`endif
